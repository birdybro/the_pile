  library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;
 
  package huffman_types is 

  type slen_type1 is array (0 to 1,0 to 15) of integer;
  constant slen : slen_type1 := ((0,0,0,0,3,1,1,1,2,2,2,3,3,3,4,4),
                                 (0,1,2,3,0,1,2,3,1,2,3,1,2,3,2,3));
   
  type sfband_l_type is array(0 to 2,0 to 22) of integer;
  constant sfBandIndex_l : sfband_l_type := 
  ((0,4,8,12,16,20,24,30,36,44,52,62,74,90,110,134,162,196,238,288,342,418,576 ),
   (0,4,8,12,16,20,24,30,36,42,50,60,72,88,106,128,156,190,230,276,330,384,576 ),
   (0,4,8,12,16,20,24,30,36,44,54,66,82,102,126,156,194,240,296,364,448,550,576 ));
    
  
  type sfband_s_type is array(0 to 2,0 to 13) of integer;
  constant sfBandIndex_s : sfband_s_type :=
  ((0,4,8,12,16,22,30,40,52,66,84,106,136,192),
  (0,4,8,12,16,22,28,38,50,64,80,100,126,192),
  (0,4,8,12,16,22,30,42,58,78,104,138,180,192));

  type table_index_type is array (0 to 33,0 to 3) of integer;
  constant table : table_index_type := 
  ((0,0,0,0),(7,2,2,0),(17,3,3,0),(17,3,3,0),(0,0,0,0),
   (31,4,4,0),(31,4,4,0),(71,6,6,0),(71,6,6,0),(71,6,6,0),
   (127,8,8,0),(127,8,8,0),(127,8,8,0),(511,16,16,0),(0,0,0,0),
   (511,16,16,0),(511,16,16,1),(511,16,16,2),(511,16,16,3),(511,16,16,4),
   (511,16,16,6),(511,16,16,8),(511,16,16,10),(511,16,16,13),(512,16,16,4),
   (512,16,16,5),(512,16,16,6),(512,16,16,7),(512,16,16,8),(512,16,16,9),
   (512,16,16,11),(512,16,16,13),(31,1,16,0),(31,1,16,0));
                                        
  subtype table_type2 is std_logic_vector(7 downto 0);
  type table_type1 is array(0 to 1) of table_type2;
  
  type table1 is array (0 to 6) of table_type1;
  constant HUFFTABLE1 : table1 :=
  ((X"02",X"01"),(X"00",X"00"),(X"02",X"01"),(X"00",X"10"),(X"02",X"01"),
  (X"00",X"01"),(X"00",X"11"));
                        
  type table2 is array (0 to 16) of table_type1;
  constant HUFFTABLE2 : table2 := 
  ((X"02",X"01"),(X"00",X"00"),(X"04",X"01"),(X"02",X"01"),(X"00",X"10"),
  (X"00",X"01"),(X"02",X"01"),(X"00",X"11"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"20"),(X"00",X"21"),(X"02",X"01"),(X"00",X"12"),(X"02",X"01"),
  (X"00",X"02"),(X"00",X"22"));
 
  type table3 is array (0 to 16) of table_type1;
  constant HUFFTABLE3 : table3 := 
  ((X"04",X"01"),(X"02",X"01"),(X"00",X"00"),(X"00",X"01"),(X"02",X"01"),
  (X"00",X"11"),(X"02",X"01"),(X"00",X"10"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"20"),(X"00",X"21"),(X"02",X"01"),(X"00",X"12"),(X"02",X"01"),
  (X"00",X"02"),(X"00",X"22"));
  
  type table5 is array (0 to 30) of table_type1;
  constant HUFFTABLE5 : table5 := 
  ((X"02",X"01"),(X"00",X"00"),(X"04",X"01"),(X"02",X"01"),(X"00",X"10"),
  (X"00",X"01"),(X"02",X"01"),(X"00",X"11"),(X"08",X"01"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"20"),(X"00",X"02"),(X"02",X"01"),(X"00",X"21"),
  (X"00",X"12"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"22"),
  (X"00",X"30"),(X"02",X"01"),(X"00",X"03"),(X"00",X"13"),(X"02",X"01"),
  (X"00",X"31"),(X"02",X"01"),(X"00",X"32"),(X"02",X"01"),(X"00",X"23"),
  (X"00",X"33")); 

  type table6 is array (0 to 30) of table_type1;
  constant HUFFTABLE6 : table6 := 
  ((X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"00"),(X"00",X"10"),
  (X"00",X"11"),(X"06",X"01"),(X"02",X"01"),(X"00",X"01"),(X"02",X"01"),  
  (X"00",X"20"),(X"00",X"21"),(X"06",X"01"),(X"02",X"01"),(X"00",X"12"),
  (X"02",X"01"),(X"00",X"02"),(X"00",X"22"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"31"),(X"00",X"13"),(X"04",X"01"),(X"02",X"01"),(X"00",X"30"),
  (X"00",X"32"),(X"02",X"01"),(X"00",X"23"),(X"02",X"01"),(X"00",X"03"),
  (X"00",X"33"));
 
  type table7 is array (0 to 70) of table_type1;
  constant HUFFTABLE7 : table7 := 
  ((X"02",X"01"),(X"00",X"00"),(X"04",X"01"),(X"02",X"01"),(X"00",X"10"),
  (X"00",X"01"),(X"08",X"01"),(X"02",X"01"),(X"00",X"11"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"20"),(X"00",X"02"),(X"00",X"21"),(X"12",X"01"),
  (X"06",X"01"),(X"02",X"01"),(X"00",X"12"),(X"02",X"01"),(X"00",X"22"),
  (X"00",X"30"),(X"04",X"01"),(X"02",X"01"),(X"00",X"31"),(X"00",X"13"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"03"),(X"00",X"32"),(X"02",X"01"),
  (X"00",X"23"),(X"00",X"04"),(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"40"),(X"00",X"41"),(X"02",X"01"),(X"00",X"14"),(X"02",X"01"),
  (X"00",X"42"),(X"00",X"24"),(X"0c",X"01"),(X"06",X"01"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"33"),(X"00",X"43"),(X"00",X"50"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"34"),(X"00",X"05"),(X"00",X"51"),(X"06",X"01"),
  (X"02",X"01"),(X"00",X"15"),(X"02",X"01"),(X"00",X"52"),(X"00",X"25"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"44"),(X"00",X"35"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"53"),(X"00",X"54"),(X"02",X"01"),(X"00",X"45"),
  (X"00",X"55"));
  
  type table8 is array (0 to 70) of table_type1;
  constant HUFFTABLE8 : table8 := 
  ((X"06",X"01"),(X"02",X"01"),(X"00",X"00"),(X"02",X"01"),(X"00",X"10"),
  (X"00",X"01"),(X"02",X"01"),(X"00",X"11"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"21"),(X"00",X"12"),(X"0e",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"20"),(X"00",X"02"),(X"02",X"01"),(X"00",X"22"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"30"),(X"00",X"03"),(X"02",X"01"),(X"00",X"31"),
  (X"00",X"13"),(X"0e",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"32"),(X"00",X"23"),(X"02",X"01"),(X"00",X"40"),(X"00",X"04"),
  (X"02",X"01"),(X"00",X"41"),(X"02",X"01"),(X"00",X"14"),(X"00",X"42"),
  (X"0c",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"24"),(X"02",X"01"),
  (X"00",X"33"),(X"00",X"50"),(X"04",X"01"),(X"02",X"01"),(X"00",X"43"),
  (X"00",X"34"),(X"00",X"51"),(X"06",X"01"),(X"02",X"01"),(X"00",X"15"),
  (X"02",X"01"),(X"00",X"05"),(X"00",X"52"),(X"06",X"01"),(X"02",X"01"),
  (X"00",X"25"),(X"02",X"01"),(X"00",X"44"),(X"00",X"35"),(X"02",X"01"),
  (X"00",X"53"),(X"02",X"01"),(X"00",X"45"),(X"02",X"01"),(X"00",X"54"),
  (X"00",X"55")); 

  type table9 is array (0 to 70) of table_type1;
  constant HUFFTABLE9 : table9 := 
  ((X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"00"),(X"00",X"10"),
(X"02",X"01"),(X"00",X"01"),(X"00",X"11"),(X"0a",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"20"),(X"00",X"21"),(X"02",X"01"),(X"00",X"12"),
(X"02",X"01"),(X"00",X"02"),(X"00",X"22"),(X"0c",X"01"),(X"06",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"30"),(X"00",X"03"),(X"00",X"31"),
(X"02",X"01"),(X"00",X"13"),(X"02",X"01"),(X"00",X"32"),(X"00",X"23"),
(X"0c",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"41"),(X"00",X"14"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"40"),(X"00",X"33"),(X"02",X"01"),
(X"00",X"42"),(X"00",X"24"),(X"0a",X"01"),(X"06",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"04"),(X"00",X"50"),(X"00",X"43"),(X"02",X"01"),
(X"00",X"34"),(X"00",X"51"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"15"),(X"00",X"52"),(X"02",X"01"),(X"00",X"25"),(X"00",X"44"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"05"),(X"00",X"54"),
(X"00",X"53"),(X"02",X"01"),(X"00",X"35"),(X"02",X"01"),(X"00",X"45"),
(X"00",X"55"));
  
  type table10 is array (0 to 126) of table_type1;
  constant HUFFTABLE10 : table10 := 
  ((X"02",X"01"),(X"00",X"00"),(X"04",X"01"),(X"02",X"01"),(X"00",X"10"),
(X"00",X"01"),(X"0a",X"01"),(X"02",X"01"),(X"00",X"11"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"20"),(X"00",X"02"),(X"02",X"01"),(X"00",X"21"),
(X"00",X"12"),(X"1c",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"22"),(X"00",X"30"),(X"02",X"01"),(X"00",X"31"),(X"00",X"13"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"03"),(X"00",X"32"),
(X"02",X"01"),(X"00",X"23"),(X"00",X"40"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"41"),(X"00",X"14"),(X"04",X"01"),(X"02",X"01"),(X"00",X"04"),
(X"00",X"33"),(X"02",X"01"),(X"00",X"42"),(X"00",X"24"),(X"1c",X"01"),
(X"0a",X"01"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"50"),
(X"00",X"05"),(X"00",X"60"),(X"02",X"01"),(X"00",X"61"),(X"00",X"16"),
(X"0c",X"01"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"43"),
(X"00",X"34"),(X"00",X"51"),(X"02",X"01"),(X"00",X"15"),(X"02",X"01"),
(X"00",X"52"),(X"00",X"25"),(X"04",X"01"),(X"02",X"01"),(X"00",X"26"),
(X"00",X"36"),(X"00",X"71"),(X"14",X"01"),(X"08",X"01"),(X"02",X"01"),
(X"00",X"17"),(X"04",X"01"),(X"02",X"01"),(X"00",X"44"),(X"00",X"53"),
(X"00",X"06"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"35"),
(X"00",X"45"),(X"00",X"62"),(X"02",X"01"),(X"00",X"70"),(X"02",X"01"),
(X"00",X"07"),(X"00",X"64"),(X"0e",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"72"),(X"00",X"27"),(X"06",X"01"),(X"02",X"01"),(X"00",X"63"),
(X"02",X"01"),(X"00",X"54"),(X"00",X"55"),(X"02",X"01"),(X"00",X"46"),
(X"00",X"73"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"37"),
(X"00",X"65"),(X"02",X"01"),(X"00",X"56"),(X"00",X"74"),(X"06",X"01"),
(X"02",X"01"),(X"00",X"47"),(X"02",X"01"),(X"00",X"66"),(X"00",X"75"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"57"),(X"00",X"76"),(X"02",X"01"),
(X"00",X"67"),(X"00",X"77")); 

  type table11 is array (0 to 126) of table_type1;
  constant HUFFTABLE11 : table11 := 
  ((X"06",X"01"),(X"02",X"01"),(X"00",X"00"),(X"02",X"01"),(X"00",X"10"),
(X"00",X"01"),(X"08",X"01"),(X"02",X"01"),(X"00",X"11"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"20"),(X"00",X"02"),(X"00",X"12"),(X"18",X"01"),
(X"08",X"01"),(X"02",X"01"),(X"00",X"21"),(X"02",X"01"),(X"00",X"22"),
(X"02",X"01"),(X"00",X"30"),(X"00",X"03"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"31"),(X"00",X"13"),(X"04",X"01"),(X"02",X"01"),(X"00",X"32"),
(X"00",X"23"),(X"04",X"01"),(X"02",X"01"),(X"00",X"40"),(X"00",X"04"),
(X"02",X"01"),(X"00",X"41"),(X"00",X"14"),(X"1e",X"01"),(X"10",X"01"),
(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"42"),(X"00",X"24"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"33"),(X"00",X"43"),(X"00",X"50"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"34"),(X"00",X"51"),(X"00",X"61"),
(X"06",X"01"),(X"02",X"01"),(X"00",X"16"),(X"02",X"01"),(X"00",X"06"),
(X"00",X"26"),(X"02",X"01"),(X"00",X"62"),(X"02",X"01"),(X"00",X"15"),
(X"02",X"01"),(X"00",X"05"),(X"00",X"52"),(X"10",X"01"),(X"0a",X"01"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"25"),(X"00",X"44"),
(X"00",X"60"),(X"02",X"01"),(X"00",X"63"),(X"00",X"36"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"70"),(X"00",X"17"),(X"00",X"71"),(X"10",X"01"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"07"),(X"00",X"64"),
(X"00",X"72"),(X"02",X"01"),(X"00",X"27"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"53"),(X"00",X"35"),(X"02",X"01"),(X"00",X"54"),(X"00",X"45"),
(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"46"),(X"00",X"73"),
(X"02",X"01"),(X"00",X"37"),(X"02",X"01"),(X"00",X"65"),(X"00",X"56"),
(X"0a",X"01"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"55"),
(X"00",X"57"),(X"00",X"74"),(X"02",X"01"),(X"00",X"47"),(X"00",X"66"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"75"),(X"00",X"76"),(X"02",X"01"),
(X"00",X"67"),(X"00",X"77"));
  
  type table12 is array (0 to 126) of table_type1;
  constant HUFFTABLE12 : table12 := 
  ((X"0c",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"10"),(X"00",X"01"),
(X"02",X"01"),(X"00",X"11"),(X"02",X"01"),(X"00",X"00"),(X"02",X"01"),
(X"00",X"20"),(X"00",X"02"),(X"10",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"21"),(X"00",X"12"),(X"04",X"01"),(X"02",X"01"),(X"00",X"22"),
(X"00",X"31"),(X"02",X"01"),(X"00",X"13"),(X"02",X"01"),(X"00",X"30"),
(X"02",X"01"),(X"00",X"03"),(X"00",X"40"),(X"1a",X"01"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"32"),(X"00",X"23"),(X"02",X"01"),
(X"00",X"41"),(X"00",X"33"),(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"14"),(X"00",X"42"),(X"02",X"01"),(X"00",X"24"),(X"02",X"01"),
(X"00",X"04"),(X"00",X"50"),(X"04",X"01"),(X"02",X"01"),(X"00",X"43"),
(X"00",X"34"),(X"02",X"01"),(X"00",X"51"),(X"00",X"15"),(X"1c",X"01"),
(X"0e",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"52"),
(X"00",X"25"),(X"02",X"01"),(X"00",X"53"),(X"00",X"35"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"60"),(X"00",X"16"),(X"00",X"61"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"62"),(X"00",X"26"),(X"06",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"05"),(X"00",X"06"),(X"00",X"44"),(X"02",X"01"),
(X"00",X"54"),(X"00",X"45"),(X"12",X"01"),(X"0a",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"63"),(X"00",X"36"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"70"),(X"00",X"07"),(X"00",X"71"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"17"),(X"00",X"64"),(X"02",X"01"),(X"00",X"46"),(X"00",X"72"),
(X"0a",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"27"),(X"02",X"01"),
(X"00",X"55"),(X"00",X"73"),(X"02",X"01"),(X"00",X"37"),(X"00",X"56"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"65"),(X"00",X"74"),
(X"02",X"01"),(X"00",X"47"),(X"00",X"66"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"75"),(X"00",X"57"),(X"02",X"01"),(X"00",X"76"),(X"02",X"01"),
(X"00",X"67"),(X"00",X"77"));

  type table13 is array (0 to 510) of table_type1;
  constant HUFFTABLE13 : table13 := 
  ((X"02",X"01"),(X"00",X"00"),(X"06",X"01"),(X"02",X"01"),(X"00",X"10"),
(X"02",X"01"),(X"00",X"01"),(X"00",X"11"),(X"1c",X"01"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"20"),(X"00",X"02"),(X"02",X"01"),
(X"00",X"21"),(X"00",X"12"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"22"),(X"00",X"30"),(X"02",X"01"),(X"00",X"03"),(X"00",X"31"),
(X"06",X"01"),(X"02",X"01"),(X"00",X"13"),(X"02",X"01"),(X"00",X"32"),
(X"00",X"23"),(X"04",X"01"),(X"02",X"01"),(X"00",X"40"),(X"00",X"04"),
(X"00",X"41"),(X"46",X"01"),(X"1c",X"01"),(X"0e",X"01"),(X"06",X"01"),
(X"02",X"01"),(X"00",X"14"),(X"02",X"01"),(X"00",X"33"),(X"00",X"42"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"24"),(X"00",X"50"),(X"02",X"01"),
(X"00",X"43"),(X"00",X"34"),(X"04",X"01"),(X"02",X"01"),(X"00",X"51"),
(X"00",X"15"),(X"04",X"01"),(X"02",X"01"),(X"00",X"05"),(X"00",X"52"),
(X"02",X"01"),(X"00",X"25"),(X"02",X"01"),(X"00",X"44"),(X"00",X"53"),
(X"0e",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"60"),
(X"00",X"06"),(X"02",X"01"),(X"00",X"61"),(X"00",X"16"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"80"),(X"00",X"08"),(X"00",X"81"),(X"10",X"01"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"35"),(X"00",X"62"),
(X"02",X"01"),(X"00",X"26"),(X"00",X"54"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"45"),(X"00",X"63"),(X"02",X"01"),(X"00",X"36"),(X"00",X"70"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"07"),(X"00",X"55"),
(X"00",X"71"),(X"02",X"01"),(X"00",X"17"),(X"02",X"01"),(X"00",X"27"),
(X"00",X"37"),(X"48",X"01"),(X"18",X"01"),(X"0c",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"18"),(X"00",X"82"),(X"02",X"01"),(X"00",X"28"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"64"),(X"00",X"46"),(X"00",X"72"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"84"),(X"00",X"48"),
(X"02",X"01"),(X"00",X"90"),(X"00",X"09"),(X"02",X"01"),(X"00",X"91"),
(X"00",X"19"),(X"18",X"01"),(X"0e",X"01"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"73"),(X"00",X"65"),(X"02",X"01"),(X"00",X"56"),
(X"00",X"74"),(X"04",X"01"),(X"02",X"01"),(X"00",X"47"),(X"00",X"66"),
(X"00",X"83"),(X"06",X"01"),(X"02",X"01"),(X"00",X"38"),(X"02",X"01"),
(X"00",X"75"),(X"00",X"57"),(X"02",X"01"),(X"00",X"92"),(X"00",X"29"),
(X"0e",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"67"),
(X"00",X"85"),(X"02",X"01"),(X"00",X"58"),(X"00",X"39"),(X"02",X"01"),
(X"00",X"93"),(X"02",X"01"),(X"00",X"49"),(X"00",X"86"),(X"06",X"01"),
(X"02",X"01"),(X"00",X"a0"),(X"02",X"01"),(X"00",X"68"),(X"00",X"0a"),
(X"02",X"01"),(X"00",X"a1"),(X"00",X"1a"),(X"44",X"01"),(X"18",X"01"),
(X"0c",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"a2"),(X"00",X"2a"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"95"),(X"00",X"59"),(X"02",X"01"),
(X"00",X"a3"),(X"00",X"3a"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"4a"),(X"00",X"96"),(X"02",X"01"),(X"00",X"b0"),(X"00",X"0b"),
(X"02",X"01"),(X"00",X"b1"),(X"00",X"1b"),(X"14",X"01"),(X"08",X"01"),
(X"02",X"01"),(X"00",X"b2"),(X"04",X"01"),(X"02",X"01"),(X"00",X"76"),
(X"00",X"77"),(X"00",X"94"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"87"),(X"00",X"78"),(X"00",X"a4"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"69"),(X"00",X"a5"),(X"00",X"2b"),(X"0c",X"01"),(X"06",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"5a"),(X"00",X"88"),(X"00",X"b3"),
(X"02",X"01"),(X"00",X"3b"),(X"02",X"01"),(X"00",X"79"),(X"00",X"a6"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"6a"),(X"00",X"b4"),
(X"00",X"c0"),(X"04",X"01"),(X"02",X"01"),(X"00",X"0c"),(X"00",X"98"),
(X"00",X"c1"),(X"3c",X"01"),(X"16",X"01"),(X"0a",X"01"),(X"06",X"01"),
(X"02",X"01"),(X"00",X"1c"),(X"02",X"01"),(X"00",X"89"),(X"00",X"b5"),
(X"02",X"01"),(X"00",X"5b"),(X"00",X"c2"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"2c"),(X"00",X"3c"),(X"04",X"01"),(X"02",X"01"),(X"00",X"b6"),
(X"00",X"6b"),(X"02",X"01"),(X"00",X"c4"),(X"00",X"4c"),(X"10",X"01"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"a8"),(X"00",X"8a"),
(X"02",X"01"),(X"00",X"d0"),(X"00",X"0d"),(X"02",X"01"),(X"00",X"d1"),
(X"02",X"01"),(X"00",X"4b"),(X"02",X"01"),(X"00",X"97"),(X"00",X"a7"),
(X"0c",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"c3"),(X"02",X"01"),
(X"00",X"7a"),(X"00",X"99"),(X"04",X"01"),(X"02",X"01"),(X"00",X"c5"),
(X"00",X"5c"),(X"00",X"b7"),(X"04",X"01"),(X"02",X"01"),(X"00",X"1d"),
(X"00",X"d2"),(X"02",X"01"),(X"00",X"2d"),(X"02",X"01"),(X"00",X"7b"),
(X"00",X"d3"),(X"34",X"01"),(X"1c",X"01"),(X"0c",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"3d"),(X"00",X"c6"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"6c"),(X"00",X"a9"),(X"02",X"01"),(X"00",X"9a"),(X"00",X"d4"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"b8"),(X"00",X"8b"),
(X"02",X"01"),(X"00",X"4d"),(X"00",X"c7"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"7c"),(X"00",X"d5"),(X"02",X"01"),(X"00",X"5d"),(X"00",X"e0"),
(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"e1"),(X"00",X"1e"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"0e"),(X"00",X"2e"),(X"00",X"e2"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"e3"),(X"00",X"6d"),
(X"02",X"01"),(X"00",X"8c"),(X"00",X"e4"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"e5"),(X"00",X"ba"),(X"00",X"f0"),(X"26",X"01"),(X"10",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"f1"),(X"00",X"1f"),(X"06",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"aa"),(X"00",X"9b"),(X"00",X"b9"),
(X"02",X"01"),(X"00",X"3e"),(X"02",X"01"),(X"00",X"d6"),(X"00",X"c8"),
(X"0c",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"4e"),(X"02",X"01"),
(X"00",X"d7"),(X"00",X"7d"),(X"02",X"01"),(X"00",X"ab"),(X"02",X"01"),
(X"00",X"5e"),(X"00",X"c9"),(X"06",X"01"),(X"02",X"01"),(X"00",X"0f"),
(X"02",X"01"),(X"00",X"9c"),(X"00",X"6e"),(X"02",X"01"),(X"00",X"f2"),
(X"00",X"2f"),(X"20",X"01"),(X"10",X"01"),(X"06",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"d8"),(X"00",X"8d"),(X"00",X"3f"),(X"06",X"01"),
(X"02",X"01"),(X"00",X"f3"),(X"02",X"01"),(X"00",X"e6"),(X"00",X"ca"),
(X"02",X"01"),(X"00",X"f4"),(X"00",X"4f"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"bb"),(X"00",X"ac"),(X"02",X"01"),(X"00",X"e7"),
(X"00",X"f5"),(X"04",X"01"),(X"02",X"01"),(X"00",X"d9"),(X"00",X"9d"),
(X"02",X"01"),(X"00",X"5f"),(X"00",X"e8"),(X"1e",X"01"),(X"0c",X"01"),
(X"06",X"01"),(X"02",X"01"),(X"00",X"6f"),(X"02",X"01"),(X"00",X"f6"),
(X"00",X"cb"),(X"04",X"01"),(X"02",X"01"),(X"00",X"bc"),(X"00",X"ad"),
(X"00",X"da"),(X"08",X"01"),(X"02",X"01"),(X"00",X"f7"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"7e"),(X"00",X"7f"),(X"00",X"8e"),(X"06",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"9e"),(X"00",X"ae"),(X"00",X"cc"),
(X"02",X"01"),(X"00",X"f8"),(X"00",X"8f"),(X"12",X"01"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"db"),(X"00",X"bd"),(X"02",X"01"),
(X"00",X"ea"),(X"00",X"f9"),(X"04",X"01"),(X"02",X"01"),(X"00",X"9f"),
(X"00",X"eb"),(X"02",X"01"),(X"00",X"be"),(X"02",X"01"),(X"00",X"cd"),
(X"00",X"fa"),(X"0e",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"dd"),
(X"00",X"ec"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"e9"),
(X"00",X"af"),(X"00",X"dc"),(X"02",X"01"),(X"00",X"ce"),(X"00",X"fb"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"bf"),(X"00",X"de"),
(X"02",X"01"),(X"00",X"cf"),(X"00",X"ee"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"df"),(X"00",X"ef"),(X"02",X"01"),(X"00",X"ff"),(X"02",X"01"),
(X"00",X"ed"),(X"02",X"01"),(X"00",X"fd"),(X"02",X"01"),(X"00",X"fc"),
(X"00",X"fe"));

  type table15 is array (0 to 510) of table_type1;
  constant HUFFTABLE15 : table15 := 
  ((X"10",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"00"),(X"02",X"01"),
(X"00",X"10"),(X"00",X"01"),(X"02",X"01"),(X"00",X"11"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"20"),(X"00",X"02"),(X"02",X"01"),(X"00",X"21"),
(X"00",X"12"),(X"32",X"01"),(X"10",X"01"),(X"06",X"01"),(X"02",X"01"),
(X"00",X"22"),(X"02",X"01"),(X"00",X"30"),(X"00",X"31"),(X"06",X"01"),
(X"02",X"01"),(X"00",X"13"),(X"02",X"01"),(X"00",X"03"),(X"00",X"40"),
(X"02",X"01"),(X"00",X"32"),(X"00",X"23"),(X"0e",X"01"),(X"06",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"04"),(X"00",X"14"),(X"00",X"41"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"33"),(X"00",X"42"),(X"02",X"01"),
(X"00",X"24"),(X"00",X"43"),(X"0a",X"01"),(X"06",X"01"),(X"02",X"01"),
(X"00",X"34"),(X"02",X"01"),(X"00",X"50"),(X"00",X"05"),(X"02",X"01"),
(X"00",X"51"),(X"00",X"15"),(X"04",X"01"),(X"02",X"01"),(X"00",X"52"),
(X"00",X"25"),(X"04",X"01"),(X"02",X"01"),(X"00",X"44"),(X"00",X"53"),
(X"00",X"61"),(X"5a",X"01"),(X"24",X"01"),(X"12",X"01"),(X"0a",X"01"),
(X"06",X"01"),(X"02",X"01"),(X"00",X"35"),(X"02",X"01"),(X"00",X"60"),
(X"00",X"06"),(X"02",X"01"),(X"00",X"16"),(X"00",X"62"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"26"),(X"00",X"54"),(X"02",X"01"),(X"00",X"45"),
(X"00",X"63"),(X"0a",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"36"),
(X"02",X"01"),(X"00",X"70"),(X"00",X"07"),(X"02",X"01"),(X"00",X"71"),
(X"00",X"55"),(X"04",X"01"),(X"02",X"01"),(X"00",X"17"),(X"00",X"64"),
(X"02",X"01"),(X"00",X"72"),(X"00",X"27"),(X"18",X"01"),(X"10",X"01"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"46"),(X"00",X"73"),
(X"02",X"01"),(X"00",X"37"),(X"00",X"65"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"56"),(X"00",X"80"),(X"02",X"01"),(X"00",X"08"),(X"00",X"74"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"81"),(X"00",X"18"),(X"02",X"01"),
(X"00",X"82"),(X"00",X"28"),(X"10",X"01"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"47"),(X"00",X"66"),(X"02",X"01"),(X"00",X"83"),
(X"00",X"38"),(X"04",X"01"),(X"02",X"01"),(X"00",X"75"),(X"00",X"57"),
(X"02",X"01"),(X"00",X"84"),(X"00",X"48"),(X"06",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"90"),(X"00",X"19"),(X"00",X"91"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"92"),(X"00",X"76"),(X"02",X"01"),(X"00",X"67"),
(X"00",X"29"),(X"5c",X"01"),(X"24",X"01"),(X"12",X"01"),(X"0a",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"85"),(X"00",X"58"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"09"),(X"00",X"77"),(X"00",X"93"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"39"),(X"00",X"94"),(X"02",X"01"),(X"00",X"49"),
(X"00",X"86"),(X"0a",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"68"),
(X"02",X"01"),(X"00",X"a0"),(X"00",X"0a"),(X"02",X"01"),(X"00",X"a1"),
(X"00",X"1a"),(X"04",X"01"),(X"02",X"01"),(X"00",X"a2"),(X"00",X"2a"),
(X"02",X"01"),(X"00",X"95"),(X"00",X"59"),(X"1a",X"01"),(X"0e",X"01"),
(X"06",X"01"),(X"02",X"01"),(X"00",X"a3"),(X"02",X"01"),(X"00",X"3a"),
(X"00",X"87"),(X"04",X"01"),(X"02",X"01"),(X"00",X"78"),(X"00",X"a4"),
(X"02",X"01"),(X"00",X"4a"),(X"00",X"96"),(X"06",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"69"),(X"00",X"b0"),(X"00",X"b1"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"1b"),(X"00",X"a5"),(X"00",X"b2"),(X"0e",X"01"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"5a"),(X"00",X"2b"),
(X"02",X"01"),(X"00",X"88"),(X"00",X"97"),(X"02",X"01"),(X"00",X"b3"),
(X"02",X"01"),(X"00",X"79"),(X"00",X"3b"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"6a"),(X"00",X"b4"),(X"02",X"01"),(X"00",X"4b"),
(X"00",X"c1"),(X"04",X"01"),(X"02",X"01"),(X"00",X"98"),(X"00",X"89"),
(X"02",X"01"),(X"00",X"1c"),(X"00",X"b5"),(X"50",X"01"),(X"22",X"01"),
(X"10",X"01"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"5b"),
(X"00",X"2c"),(X"00",X"c2"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"0b"),(X"00",X"c0"),(X"00",X"a6"),(X"02",X"01"),(X"00",X"a7"),
(X"00",X"7a"),(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"c3"),
(X"00",X"3c"),(X"04",X"01"),(X"02",X"01"),(X"00",X"0c"),(X"00",X"99"),
(X"00",X"b6"),(X"04",X"01"),(X"02",X"01"),(X"00",X"6b"),(X"00",X"c4"),
(X"02",X"01"),(X"00",X"4c"),(X"00",X"a8"),(X"14",X"01"),(X"0a",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"8a"),(X"00",X"c5"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"d0"),(X"00",X"5c"),(X"00",X"d1"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"b7"),(X"00",X"7b"),(X"02",X"01"),(X"00",X"1d"),
(X"02",X"01"),(X"00",X"0d"),(X"00",X"2d"),(X"0c",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"d2"),(X"00",X"d3"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"3d"),(X"00",X"c6"),(X"02",X"01"),(X"00",X"6c"),(X"00",X"a9"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"9a"),(X"00",X"b8"),
(X"00",X"d4"),(X"04",X"01"),(X"02",X"01"),(X"00",X"8b"),(X"00",X"4d"),
(X"02",X"01"),(X"00",X"c7"),(X"00",X"7c"),(X"44",X"01"),(X"22",X"01"),
(X"12",X"01"),(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"d5"),
(X"00",X"5d"),(X"04",X"01"),(X"02",X"01"),(X"00",X"e0"),(X"00",X"0e"),
(X"00",X"e1"),(X"04",X"01"),(X"02",X"01"),(X"00",X"1e"),(X"00",X"e2"),
(X"02",X"01"),(X"00",X"aa"),(X"00",X"2e"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"b9"),(X"00",X"9b"),(X"02",X"01"),(X"00",X"e3"),
(X"00",X"d6"),(X"04",X"01"),(X"02",X"01"),(X"00",X"6d"),(X"00",X"3e"),
(X"02",X"01"),(X"00",X"c8"),(X"00",X"8c"),(X"10",X"01"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"e4"),(X"00",X"4e"),(X"02",X"01"),
(X"00",X"d7"),(X"00",X"7d"),(X"04",X"01"),(X"02",X"01"),(X"00",X"e5"),
(X"00",X"ba"),(X"02",X"01"),(X"00",X"ab"),(X"00",X"5e"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"c9"),(X"00",X"9c"),(X"02",X"01"),
(X"00",X"f1"),(X"00",X"1f"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"f0"),(X"00",X"6e"),(X"00",X"f2"),(X"02",X"01"),(X"00",X"2f"),
(X"00",X"e6"),(X"26",X"01"),(X"12",X"01"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"d8"),(X"00",X"f3"),(X"02",X"01"),(X"00",X"3f"),
(X"00",X"f4"),(X"06",X"01"),(X"02",X"01"),(X"00",X"4f"),(X"02",X"01"),
(X"00",X"8d"),(X"00",X"d9"),(X"02",X"01"),(X"00",X"bb"),(X"00",X"ca"),
(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"ac"),(X"00",X"e7"),
(X"02",X"01"),(X"00",X"7e"),(X"00",X"f5"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"9d"),(X"00",X"5f"),(X"02",X"01"),(X"00",X"e8"),
(X"00",X"8e"),(X"02",X"01"),(X"00",X"f6"),(X"00",X"cb"),(X"22",X"01"),
(X"12",X"01"),(X"0a",X"01"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"0f"),(X"00",X"ae"),(X"00",X"6f"),(X"02",X"01"),(X"00",X"bc"),
(X"00",X"da"),(X"04",X"01"),(X"02",X"01"),(X"00",X"ad"),(X"00",X"f7"),
(X"02",X"01"),(X"00",X"7f"),(X"00",X"e9"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"9e"),(X"00",X"cc"),(X"02",X"01"),(X"00",X"f8"),
(X"00",X"8f"),(X"04",X"01"),(X"02",X"01"),(X"00",X"db"),(X"00",X"bd"),
(X"02",X"01"),(X"00",X"ea"),(X"00",X"f9"),(X"10",X"01"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"9f"),(X"00",X"dc"),(X"02",X"01"),
(X"00",X"cd"),(X"00",X"eb"),(X"04",X"01"),(X"02",X"01"),(X"00",X"be"),
(X"00",X"fa"),(X"02",X"01"),(X"00",X"af"),(X"00",X"dd"),(X"0e",X"01"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"ec"),(X"00",X"ce"),
(X"00",X"fb"),(X"04",X"01"),(X"02",X"01"),(X"00",X"bf"),(X"00",X"ed"),
(X"02",X"01"),(X"00",X"de"),(X"00",X"fc"),(X"06",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"cf"),(X"00",X"fd"),(X"00",X"ee"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"df"),(X"00",X"fe"),(X"02",X"01"),(X"00",X"ef"),
(X"00",X"ff"));
  
  type table16 is array (0 to 510) of table_type1;
  constant HUFFTABLE16 : table16 := 
  ((X"02",X"01"),(X"00",X"00"),(X"06",X"01"),(X"02",X"01"),(X"00",X"10"),
(X"02",X"01"),(X"00",X"01"),(X"00",X"11"),(X"2a",X"01"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"20"),(X"00",X"02"),(X"02",X"01"),
(X"00",X"21"),(X"00",X"12"),(X"0a",X"01"),(X"06",X"01"),(X"02",X"01"),
(X"00",X"22"),(X"02",X"01"),(X"00",X"30"),(X"00",X"03"),(X"02",X"01"),
(X"00",X"31"),(X"00",X"13"),(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"32"),(X"00",X"23"),(X"04",X"01"),(X"02",X"01"),(X"00",X"40"),
(X"00",X"04"),(X"00",X"41"),(X"06",X"01"),(X"02",X"01"),(X"00",X"14"),
(X"02",X"01"),(X"00",X"33"),(X"00",X"42"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"24"),(X"00",X"50"),(X"02",X"01"),(X"00",X"43"),(X"00",X"34"),
(X"8a",X"01"),(X"28",X"01"),(X"10",X"01"),(X"06",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"05"),(X"00",X"15"),(X"00",X"51"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"52"),(X"00",X"25"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"44"),(X"00",X"35"),(X"00",X"53"),(X"0a",X"01"),(X"06",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"60"),(X"00",X"06"),(X"00",X"61"),
(X"02",X"01"),(X"00",X"16"),(X"00",X"62"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"26"),(X"00",X"54"),(X"02",X"01"),(X"00",X"45"),
(X"00",X"63"),(X"04",X"01"),(X"02",X"01"),(X"00",X"36"),(X"00",X"70"),
(X"00",X"71"),(X"28",X"01"),(X"12",X"01"),(X"08",X"01"),(X"02",X"01"),
(X"00",X"17"),(X"02",X"01"),(X"00",X"07"),(X"02",X"01"),(X"00",X"55"),
(X"00",X"64"),(X"04",X"01"),(X"02",X"01"),(X"00",X"72"),(X"00",X"27"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"46"),(X"00",X"65"),(X"00",X"73"),
(X"0a",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"37"),(X"02",X"01"),
(X"00",X"56"),(X"00",X"08"),(X"02",X"01"),(X"00",X"80"),(X"00",X"81"),
(X"06",X"01"),(X"02",X"01"),(X"00",X"18"),(X"02",X"01"),(X"00",X"74"),
(X"00",X"47"),(X"02",X"01"),(X"00",X"82"),(X"02",X"01"),(X"00",X"28"),
(X"00",X"66"),(X"18",X"01"),(X"0e",X"01"),(X"08",X"01"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"83"),(X"00",X"38"),(X"02",X"01"),(X"00",X"75"),
(X"00",X"84"),(X"04",X"01"),(X"02",X"01"),(X"00",X"48"),(X"00",X"90"),
(X"00",X"91"),(X"06",X"01"),(X"02",X"01"),(X"00",X"19"),(X"02",X"01"),
(X"00",X"09"),(X"00",X"76"),(X"02",X"01"),(X"00",X"92"),(X"00",X"29"),
(X"0e",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"85"),
(X"00",X"58"),(X"02",X"01"),(X"00",X"93"),(X"00",X"39"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"a0"),(X"00",X"0a"),(X"00",X"1a"),(X"08",X"01"),
(X"02",X"01"),(X"00",X"a2"),(X"02",X"01"),(X"00",X"67"),(X"02",X"01"),
(X"00",X"57"),(X"00",X"49"),(X"06",X"01"),(X"02",X"01"),(X"00",X"94"),
(X"02",X"01"),(X"00",X"77"),(X"00",X"86"),(X"02",X"01"),(X"00",X"a1"),
(X"02",X"01"),(X"00",X"68"),(X"00",X"95"),(X"dc",X"01"),(X"7e",X"01"),
(X"32",X"01"),(X"1a",X"01"),(X"0c",X"01"),(X"06",X"01"),(X"02",X"01"),
(X"00",X"2a"),(X"02",X"01"),(X"00",X"59"),(X"00",X"3a"),(X"02",X"01"),
(X"00",X"a3"),(X"02",X"01"),(X"00",X"87"),(X"00",X"78"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"a4"),(X"00",X"4a"),(X"02",X"01"),
(X"00",X"96"),(X"00",X"69"),(X"04",X"01"),(X"02",X"01"),(X"00",X"b0"),
(X"00",X"0b"),(X"00",X"b1"),(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"1b"),(X"00",X"b2"),(X"02",X"01"),(X"00",X"2b"),(X"02",X"01"),
(X"00",X"a5"),(X"00",X"5a"),(X"06",X"01"),(X"02",X"01"),(X"00",X"b3"),
(X"02",X"01"),(X"00",X"a6"),(X"00",X"6a"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"b4"),(X"00",X"4b"),(X"02",X"01"),(X"00",X"0c"),(X"00",X"c1"),
(X"1e",X"01"),(X"0e",X"01"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"b5"),(X"00",X"c2"),(X"00",X"2c"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"a7"),(X"00",X"c3"),(X"02",X"01"),(X"00",X"6b"),(X"00",X"c4"),
(X"08",X"01"),(X"02",X"01"),(X"00",X"1d"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"88"),(X"00",X"97"),(X"00",X"3b"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"d1"),(X"00",X"d2"),(X"02",X"01"),(X"00",X"2d"),(X"00",X"d3"),
(X"12",X"01"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"1e"),
(X"00",X"2e"),(X"00",X"e2"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"79"),(X"00",X"98"),(X"00",X"c0"),(X"02",X"01"),(X"00",X"1c"),
(X"02",X"01"),(X"00",X"89"),(X"00",X"5b"),(X"0e",X"01"),(X"06",X"01"),
(X"02",X"01"),(X"00",X"3c"),(X"02",X"01"),(X"00",X"7a"),(X"00",X"b6"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"4c"),(X"00",X"99"),(X"02",X"01"),
(X"00",X"a8"),(X"00",X"8a"),(X"06",X"01"),(X"02",X"01"),(X"00",X"0d"),
(X"02",X"01"),(X"00",X"c5"),(X"00",X"5c"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"3d"),(X"00",X"c6"),(X"02",X"01"),(X"00",X"6c"),(X"00",X"9a"),
(X"58",X"01"),(X"56",X"01"),(X"24",X"01"),(X"10",X"01"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"8b"),(X"00",X"4d"),(X"02",X"01"),
(X"00",X"c7"),(X"00",X"7c"),(X"04",X"01"),(X"02",X"01"),(X"00",X"d5"),
(X"00",X"5d"),(X"02",X"01"),(X"00",X"e0"),(X"00",X"0e"),(X"08",X"01"),
(X"02",X"01"),(X"00",X"e3"),(X"04",X"01"),(X"02",X"01"),(X"00",X"d0"),
(X"00",X"b7"),(X"00",X"7b"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"a9"),(X"00",X"b8"),(X"00",X"d4"),(X"02",X"01"),(X"00",X"e1"),
(X"02",X"01"),(X"00",X"aa"),(X"00",X"b9"),(X"18",X"01"),(X"0a",X"01"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"9b"),(X"00",X"d6"),
(X"00",X"6d"),(X"02",X"01"),(X"00",X"3e"),(X"00",X"c8"),(X"06",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"8c"),(X"00",X"e4"),(X"00",X"4e"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"d7"),(X"00",X"e5"),(X"02",X"01"),
(X"00",X"ba"),(X"00",X"ab"),(X"0c",X"01"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"9c"),(X"00",X"e6"),(X"04",X"01"),(X"02",X"01"),(X"00",X"6e"),
(X"00",X"d8"),(X"02",X"01"),(X"00",X"8d"),(X"00",X"bb"),(X"08",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"e7"),(X"00",X"9d"),(X"02",X"01"),
(X"00",X"e8"),(X"00",X"8e"),(X"04",X"01"),(X"02",X"01"),(X"00",X"cb"),
(X"00",X"bc"),(X"00",X"9e"),(X"00",X"f1"),(X"02",X"01"),(X"00",X"1f"),
(X"02",X"01"),(X"00",X"0f"),(X"00",X"2f"),(X"42",X"01"),(X"38",X"01"),
(X"02",X"01"),(X"00",X"f2"),(X"34",X"01"),(X"32",X"01"),(X"14",X"01"),
(X"08",X"01"),(X"02",X"01"),(X"00",X"bd"),(X"02",X"01"),(X"00",X"5e"),
(X"02",X"01"),(X"00",X"7d"),(X"00",X"c9"),(X"06",X"01"),(X"02",X"01"),
(X"00",X"ca"),(X"02",X"01"),(X"00",X"ac"),(X"00",X"7e"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"da"),(X"00",X"ad"),(X"00",X"cc"),(X"0a",X"01"),
(X"06",X"01"),(X"02",X"01"),(X"00",X"ae"),(X"02",X"01"),(X"00",X"db"),
(X"00",X"dc"),(X"02",X"01"),(X"00",X"cd"),(X"00",X"be"),(X"06",X"01"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"eb"),(X"00",X"ed"),(X"00",X"ee"),
(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"d9"),(X"00",X"ea"),
(X"00",X"e9"),(X"02",X"01"),(X"00",X"de"),(X"04",X"01"),(X"02",X"01"),
(X"00",X"dd"),(X"00",X"ec"),(X"00",X"ce"),(X"00",X"3f"),(X"00",X"f0"),
(X"04",X"01"),(X"02",X"01"),(X"00",X"f3"),(X"00",X"f4"),(X"02",X"01"),
(X"00",X"4f"),(X"02",X"01"),(X"00",X"f5"),(X"00",X"5f"),(X"0a",X"01"),
(X"02",X"01"),(X"00",X"ff"),(X"04",X"01"),(X"02",X"01"),(X"00",X"f6"),
(X"00",X"6f"),(X"02",X"01"),(X"00",X"f7"),(X"00",X"7f"),(X"0c",X"01"),
(X"06",X"01"),(X"02",X"01"),(X"00",X"8f"),(X"02",X"01"),(X"00",X"f8"),
(X"00",X"f9"),(X"04",X"01"),(X"02",X"01"),(X"00",X"9f"),(X"00",X"fa"),
(X"00",X"af"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"fb"),
(X"00",X"bf"),(X"02",X"01"),(X"00",X"fc"),(X"00",X"cf"),(X"04",X"01"),
(X"02",X"01"),(X"00",X"fd"),(X"00",X"df"),(X"02",X"01"),(X"00",X"fe"),
(X"00",X"ef"));
  
  type table24 is array (0 to 511) of table_type1;
  constant HUFFTABLE24 : table24 := 
  ((X"3c",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"00"),
  (X"00",X"10"),(X"02",X"01"),(X"00",X"01"),(X"00",X"11"),(X"0e",X"01"),
  (X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"20"),(X"00",X"02"),
  (X"00",X"21"),(X"02",X"01"),(X"00",X"12"),(X"02",X"01"),(X"00",X"22"),
  (X"02",X"01"),(X"00",X"30"),(X"00",X"03"),(X"0e",X"01"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"31"),(X"00",X"13"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"32"),(X"00",X"23"),(X"04",X"01"),(X"02",X"01"),(X"00",X"40"),
  (X"00",X"04"),(X"00",X"41"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"14"),(X"00",X"33"),(X"02",X"01"),(X"00",X"42"),(X"00",X"24"),
  (X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"43"),(X"00",X"34"),
  (X"00",X"51"),(X"06",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"50"),
  (X"00",X"05"),(X"00",X"15"),(X"02",X"01"),(X"00",X"52"),(X"00",X"25"),
  (X"fa",X"01"),(X"62",X"01"),(X"22",X"01"),(X"12",X"01"),(X"0a",X"01"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"44"),(X"00",X"53"),(X"02",X"01"),
  (X"00",X"35"),(X"02",X"01"),(X"00",X"60"),(X"00",X"06"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"61"),(X"00",X"16"),(X"02",X"01"),(X"00",X"62"),
  (X"00",X"26"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"54"),
  (X"00",X"45"),(X"02",X"01"),(X"00",X"63"),(X"00",X"36"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"71"),(X"00",X"55"),(X"02",X"01"),(X"00",X"64"),
  (X"00",X"46"),(X"20",X"01"),(X"0e",X"01"),(X"06",X"01"),(X"02",X"01"),
  (X"00",X"72"),(X"02",X"01"),(X"00",X"27"),(X"00",X"37"),(X"02",X"01"),
  (X"00",X"73"),(X"04",X"01"),(X"02",X"01"),(X"00",X"70"),(X"00",X"07"),
  (X"00",X"17"),(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"65"),
  (X"00",X"56"),(X"04",X"01"),(X"02",X"01"),(X"00",X"80"),(X"00",X"08"),
  (X"00",X"81"),(X"04",X"01"),(X"02",X"01"),(X"00",X"74"),(X"00",X"47"),
  (X"02",X"01"),(X"00",X"18"),(X"00",X"82"),(X"10",X"01"),(X"08",X"01"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"28"),(X"00",X"66"),(X"02",X"01"),
  (X"00",X"83"),(X"00",X"38"),(X"04",X"01"),(X"02",X"01"),(X"00",X"75"),
  (X"00",X"57"),(X"02",X"01"),(X"00",X"84"),(X"00",X"48"),(X"08",X"01"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"91"),(X"00",X"19"),(X"02",X"01"),
  (X"00",X"92"),(X"00",X"76"),(X"04",X"01"),(X"02",X"01"),(X"00",X"67"),
  (X"00",X"29"),(X"02",X"01"),(X"00",X"85"),(X"00",X"58"),(X"5c",X"01"),
  (X"22",X"01"),(X"10",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"93"),(X"00",X"39"),(X"02",X"01"),(X"00",X"94"),(X"00",X"49"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"77"),(X"00",X"86"),(X"02",X"01"),
  (X"00",X"68"),(X"00",X"a1"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"a2"),(X"00",X"2a"),(X"02",X"01"),(X"00",X"95"),(X"00",X"59"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"a3"),(X"00",X"3a"),(X"02",X"01"),
  (X"00",X"87"),(X"02",X"01"),(X"00",X"78"),(X"00",X"4a"),(X"16",X"01"),
  (X"0c",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"a4"),(X"00",X"96"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"69"),(X"00",X"b1"),(X"02",X"01"),
  (X"00",X"1b"),(X"00",X"a5"),(X"06",X"01"),(X"02",X"01"),(X"00",X"b2"),
  (X"02",X"01"),(X"00",X"5a"),(X"00",X"2b"),(X"02",X"01"),(X"00",X"88"),
  (X"00",X"b3"),(X"10",X"01"),(X"0a",X"01"),(X"06",X"01"),(X"02",X"01"),
  (X"00",X"90"),(X"02",X"01"),(X"00",X"09"),(X"00",X"a0"),(X"02",X"01"),
  (X"00",X"97"),(X"00",X"79"),(X"04",X"01"),(X"02",X"01"),(X"00",X"a6"),
  (X"00",X"6a"),(X"00",X"b4"),(X"0c",X"01"),(X"06",X"01"),(X"02",X"01"),
  (X"00",X"1a"),(X"02",X"01"),(X"00",X"0a"),(X"00",X"b0"),(X"02",X"01"),
  (X"00",X"3b"),(X"02",X"01"),(X"00",X"0b"),(X"00",X"c0"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"4b"),(X"00",X"c1"),(X"02",X"01"),(X"00",X"98"),
  (X"00",X"89"),(X"43",X"01"),(X"22",X"01"),(X"10",X"01"),(X"08",X"01"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"1c"),(X"00",X"b5"),(X"02",X"01"),
  (X"00",X"5b"),(X"00",X"c2"),(X"04",X"01"),(X"02",X"01"),(X"00",X"2c"),
  (X"00",X"a7"),(X"02",X"01"),(X"00",X"7a"),(X"00",X"c3"),(X"0a",X"01"),
  (X"06",X"01"),(X"02",X"01"),(X"00",X"3c"),(X"02",X"01"),(X"00",X"0c"),
  (X"00",X"d0"),(X"02",X"01"),(X"00",X"b6"),(X"00",X"6b"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"c4"),(X"00",X"4c"),(X"02",X"01"),(X"00",X"99"),
  (X"00",X"a8"),(X"10",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"8a"),(X"00",X"c5"),(X"02",X"01"),(X"00",X"5c"),(X"00",X"d1"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"b7"),(X"00",X"7b"),(X"02",X"01"),
  (X"00",X"1d"),(X"00",X"d2"),(X"09",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"2d"),(X"00",X"d3"),(X"02",X"01"),(X"00",X"3d"),(X"00",X"c6"),
  (X"55",X"fa"),(X"04",X"01"),(X"02",X"01"),(X"00",X"6c"),(X"00",X"a9"),
  (X"02",X"01"),(X"00",X"9a"),(X"00",X"d4"),(X"20",X"01"),(X"10",X"01"),
  (X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"b8"),(X"00",X"8b"),
  (X"02",X"01"),(X"00",X"4d"),(X"00",X"c7"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"7c"),(X"00",X"d5"),(X"02",X"01"),(X"00",X"5d"),(X"00",X"e1"),
  (X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"1e"),(X"00",X"e2"),
  (X"02",X"01"),(X"00",X"aa"),(X"00",X"b9"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"9b"),(X"00",X"e3"),(X"02",X"01"),(X"00",X"d6"),(X"00",X"6d"),
  (X"14",X"01"),(X"0a",X"01"),(X"06",X"01"),(X"02",X"01"),(X"00",X"3e"),
  (X"02",X"01"),(X"00",X"2e"),(X"00",X"4e"),(X"02",X"01"),(X"00",X"c8"),
  (X"00",X"8c"),(X"04",X"01"),(X"02",X"01"),(X"00",X"e4"),(X"00",X"d7"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"7d"),(X"00",X"ab"),(X"00",X"e5"),
  (X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"ba"),(X"00",X"5e"),
  (X"02",X"01"),(X"00",X"c9"),(X"02",X"01"),(X"00",X"9c"),(X"00",X"6e"),
  (X"08",X"01"),(X"02",X"01"),(X"00",X"e6"),(X"02",X"01"),(X"00",X"0d"),
  (X"02",X"01"),(X"00",X"e0"),(X"00",X"0e"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"d8"),(X"00",X"8d"),(X"02",X"01"),(X"00",X"bb"),(X"00",X"ca"),
  (X"4a",X"01"),(X"02",X"01"),(X"00",X"ff"),(X"40",X"01"),(X"3a",X"01"),
  (X"20",X"01"),(X"10",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"ac"),(X"00",X"e7"),(X"02",X"01"),(X"00",X"7e"),(X"00",X"d9"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"9d"),(X"00",X"e8"),(X"02",X"01"),
  (X"00",X"8e"),(X"00",X"cb"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"bc"),(X"00",X"da"),(X"02",X"01"),(X"00",X"ad"),(X"00",X"e9"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"9e"),(X"00",X"cc"),(X"02",X"01"),
  (X"00",X"db"),(X"00",X"bd"),(X"10",X"01"),(X"08",X"01"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"ea"),(X"00",X"ae"),(X"02",X"01"),(X"00",X"dc"),
  (X"00",X"cd"),(X"04",X"01"),(X"02",X"01"),(X"00",X"eb"),(X"00",X"be"),
  (X"02",X"01"),(X"00",X"dd"),(X"00",X"ec"),(X"08",X"01"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"ce"),(X"00",X"ed"),(X"02",X"01"),(X"00",X"de"),
  (X"00",X"ee"),(X"00",X"0f"),(X"04",X"01"),(X"02",X"01"),(X"00",X"f0"),
  (X"00",X"1f"),(X"00",X"f1"),(X"04",X"01"),(X"02",X"01"),(X"00",X"f2"),
  (X"00",X"2f"),(X"02",X"01"),(X"00",X"f3"),(X"00",X"3f"),(X"12",X"01"),
  (X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"f4"),(X"00",X"4f"),
  (X"02",X"01"),(X"00",X"f5"),(X"00",X"5f"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"f6"),(X"00",X"6f"),(X"02",X"01"),(X"00",X"f7"),(X"02",X"01"),
  (X"00",X"7f"),(X"00",X"8f"),(X"0a",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"f8"),(X"00",X"f9"),(X"04",X"01"),(X"02",X"01"),(X"00",X"9f"),
  (X"00",X"af"),(X"00",X"fa"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"fb"),(X"00",X"bf"),(X"02",X"01"),(X"00",X"fc"),(X"00",X"cf"),
  (X"04",X"01"),(X"02",X"01"),(X"00",X"fd"),(X"00",X"df"),(X"02",X"01"),
  (X"00",X"fe"),(X"00",X"ef"));

  type table32 is array (0 to 30) of table_type1;
  constant HUFFTABLE32 : table32 := 
  ((X"02",X"01"),(X"00",X"00"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),
  (X"00",X"08"),(X"00",X"04"),(X"02",X"01"),(X"00",X"01"),(X"00",X"02"),
  (X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"0c"),(X"00",X"0a"),
  (X"02",X"01"),(X"00",X"03"),(X"00",X"06"),(X"06",X"01"),(X"02",X"01"),
  (X"00",X"09"),(X"02",X"01"),(X"00",X"05"),(X"00",X"07"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"0e"),(X"00",X"0d"),(X"02",X"01"),(X"00",X"0f"),
  (X"00",X"0b"));  
 
  type table33 is array (0 to 30) of table_type1;  
  constant HUFFTABLE33 : table33 := 
  ((X"10",X"01"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"00"),
  (X"00",X"01"),(X"02",X"01"),(X"00",X"02"),(X"00",X"03"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"04"),(X"00",X"05"),(X"02",X"01"),(X"00",X"06"),
  (X"00",X"07"),(X"08",X"01"),(X"04",X"01"),(X"02",X"01"),(X"00",X"08"),
  (X"00",X"09"),(X"02",X"01"),(X"00",X"0a"),(X"00",X"0b"),(X"04",X"01"),
  (X"02",X"01"),(X"00",X"0c"),(X"00",X"0d"),(X"02",X"01"),(X"00",X"0e"),
  (X"00",X"0f"));
  
  function get_value(tindex,level,index:in integer) return integer;
end;

package body huffman_types is

function get_value(tindex,level,index:in integer) return integer is 
variable val:integer;

begin
  case tindex is 
      when 0 =>
           val :=0;     
      when 1 =>
           val := conv_integer(HUFFTABLE1(level)(index));
      when 2 => 
           val := conv_integer(HUFFTABLE2(level)(index));
      when 3 =>
           val :=conv_integer(HUFFTABLE3(level)(index));
      when 4 =>
           val :=0;
      when 5 =>
           val :=conv_integer(HUFFTABLE5(level)(index));
      when 6 =>
           val :=conv_integer(HUFFTABLE6(level)(index));
      when 7 =>
           val :=conv_integer(HUFFTABLE7(level)(index));
      when 8 =>
           val :=conv_integer(HUFFTABLE8(level)(index));
      when 9 =>
           val :=conv_integer(HUFFTABLE9(level)(index));
      when 10 =>
           val :=conv_integer(HUFFTABLE10(level)(index));
      when 11 =>
           val :=conv_integer(HUFFTABLE11(level)(index));
      when 12 =>
           val :=conv_integer(HUFFTABLE12(level)(index));
      when 13 =>
           val :=conv_integer(HUFFTABLE13(level)(index));
      when 14 =>
           val :=0;
      when 15 =>
           val :=conv_integer(HUFFTABLE15(level)(index));
      when 16 =>
           val :=conv_integer(HUFFTABLE16(level)(index));
      when 17 =>
           val :=conv_integer(HUFFTABLE16(level)(index));
      when 18 =>
           val :=conv_integer(HUFFTABLE16(level)(index));
      when 19 =>
           val :=conv_integer(HUFFTABLE16(level)(index));
      when 20 => 
           val :=conv_integer(HUFFTABLE16(level)(index));
      when 21 =>
           val :=conv_integer(HUFFTABLE16(level)(index));
      when 22 =>
           val :=conv_integer(HUFFTABLE16(level)(index));
      when 23 =>
           val :=conv_integer(HUFFTABLE16(level)(index));
      when 24 =>
           val :=conv_integer(HUFFTABLE24(level)(index));
      when 25 =>
           val :=conv_integer(HUFFTABLE24(level)(index));
      when 26 =>
           val :=conv_integer(HUFFTABLE24(level)(index));
      when 27 =>
           val :=conv_integer(HUFFTABLE24(level)(index));
      when 28 =>
           val :=conv_integer(HUFFTABLE24(level)(index));
      when 29 =>
           val :=conv_integer(HUFFTABLE24(level)(index));
      when 31 =>
           val :=conv_integer(HUFFTABLE24(level)(index));
      when 32 =>
           val :=conv_integer(HUFFTABLE32(level)(index));
      when 33 =>
           val :=conv_integer(HUFFTABLE33(level)(index));
      when others =>
    end case;

  return val;
  end function;
end package body;