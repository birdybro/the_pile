// 
//  MAC_MPEG2_AV - MPEG-2 hardware implementation for Xilinx multimedia board 
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MPEG2_AV
// 
// MAC_MPEG2_AV is distributed in the hope that it will be useful for further 
// research, but WITHOUT ANY WARRANTY; without even the implied warranty of 
//	MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. MAC_MPEG2_AV is free; you 
// can redistribute it and/or modify it provided that proper reference is provided 
// to the authors. See the documents included in the "doc" folder for further details.
//
//==============================================================================

`include "defines.v"
module Quant_Scan_ROM(
   clock,
   Enable_A_I,
   Address_A_I,
   Data_A_O,
   Enable_B_I,
   Address_B_I,
   Data_B_O
);

input             clock;
input             Enable_A_I;
input    [10:0]   Address_A_I;
output   [7:0]    Data_A_O;
input             Enable_B_I;
input    [10:0]   Address_B_I;
output   [7:0]    Data_B_O;

wire     [7:0]    Data_A, Data_B;

assign Data_A_O = Data_A;
assign Data_B_O = Data_B;

RAMB16_S9_S9 Quant_Scan_Matrix_ROM (
   .DOA(Data_A),
   .DOB(Data_B),
   .DOPA(),
   .DOPB(),
   .ADDRA(Address_A_I),
   .ADDRB(Address_B_I),
   .CLKA(clock),
   .CLKB(clock),
   .DIA(8'h00),
   .DIB(8'h00),
   .DIPA(1'b0),
   .DIPB(1'b0),
   .ENA(Enable_A_I),
   .ENB(Enable_B_I),
   .SSRA(1'b0),
   .SSRB(1'b0),
   .WEA(1'b0),
   .WEB(1'b0)
);

// synthesis attribute INIT_00 of Quant_Scan_Matrix_ROM is "256'h1C150E07060D141B22293028211A130C05040B12192018110A03020910080100"
// synthesis attribute INIT_01 of Quant_Scan_Matrix_ROM is "256'h3F3E372F363D3C352E271F262D343B3A332C251E170F161D242B323938312A23"
// synthesis attribute INIT_02 of Quant_Scan_Matrix_ROM is "256'h2B233A322A221B130C040B03121A212931393830282019110A02090118100800"
// synthesis attribute INIT_03 of Quant_Scan_Matrix_ROM is "256'h3F372F273E362E261F170F071E163D352D253C342C241D150E060D051C143B33"
// synthesis attribute INIT_04 of Quant_Scan_Matrix_ROM is "256'h2825221D1B1A16162622221D1B1A161325221D1B18161010221D1B1A16131008"
// synthesis attribute INIT_05 of Quant_Scan_Matrix_ROM is "256'h5345382E26231D1B45382E26221D1B1A3A302823201D1B1A302823201D1B1A16"
// synthesis attribute INIT_06 of Quant_Scan_Matrix_ROM is "256'h1010101010101010101010101010101010101010101010101010101010101010"
// synthesis attribute INIT_07 of Quant_Scan_Matrix_ROM is "256'h1010101010101010101010101010101010101010101010101010101010101010"
                                                                                                                                 
// synthesis attribute INIT_08 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_09 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0A of Quant_Scan_Matrix_ROM is "256'h1B19181716151413191817161514131218171615141312111716151413121110"
// synthesis attribute INIT_0B of Quant_Scan_Matrix_ROM is "256'h211F1E1C1B1918171F1E1C1B191817161E1C1B19181716151C1B191817161514"
// synthesis attribute INIT_0C of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0D of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0E of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0F of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
                                                                                                                                 
// synthesis attribute INIT_10 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_11 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_12 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_13 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_14 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_15 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_16 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_17 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
                                                                                                                                 
// synthesis attribute INIT_18 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_19 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1A of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1B of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1C of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1D of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1E of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1F of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
                                                                                                                                 
// synthesis attribute INIT_20 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_21 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_22 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_23 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_24 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_25 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_26 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_27 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
                                                                                                                                 
// synthesis attribute INIT_28 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_29 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2A of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2B of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2C of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2D of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2E of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2F of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
                                                                                                                                 
// synthesis attribute INIT_30 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_31 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_32 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_33 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_34 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_35 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_36 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_37 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
                                                                                                                                 
// synthesis attribute INIT_38 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_39 of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3A of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3B of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3C of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3D of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3E of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3F of Quant_Scan_Matrix_ROM is "256'h0000000000000000000000000000000000000000000000000000000000000000"

// synthesis translate_off

defparam Quant_Scan_Matrix_ROM.INIT_00 = 256'h1C150E07060D141B22293028211A130C05040B12192018110A03020910080100;
defparam Quant_Scan_Matrix_ROM.INIT_01 = 256'h3F3E372F363D3C352E271F262D343B3A332C251E170F161D242B323938312A23;
defparam Quant_Scan_Matrix_ROM.INIT_02 = 256'h2B233A322A221B130C040B03121A212931393830282019110A02090118100800;
defparam Quant_Scan_Matrix_ROM.INIT_03 = 256'h3F372F273E362E261F170F071E163D352D253C342C241D150E060D051C143B33;
defparam Quant_Scan_Matrix_ROM.INIT_04 = 256'h2825221D1B1A16162622221D1B1A161325221D1B18161010221D1B1A16131008;
defparam Quant_Scan_Matrix_ROM.INIT_05 = 256'h5345382E26231D1B45382E26221D1B1A3A302823201D1B1A302823201D1B1A16;
defparam Quant_Scan_Matrix_ROM.INIT_06 = 256'h1010101010101010101010101010101010101010101010101010101010101010;
defparam Quant_Scan_Matrix_ROM.INIT_07 = 256'h1010101010101010101010101010101010101010101010101010101010101010;
                                                                                                              
defparam Quant_Scan_Matrix_ROM.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_0A = 256'h1B19181716151413191817161514131218171615141312111716151413121110;
defparam Quant_Scan_Matrix_ROM.INIT_0B = 256'h211F1E1C1B1918171F1E1C1B191817161E1C1B19181716151C1B191817161514;
defparam Quant_Scan_Matrix_ROM.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                              
defparam Quant_Scan_Matrix_ROM.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                              
defparam Quant_Scan_Matrix_ROM.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                              
defparam Quant_Scan_Matrix_ROM.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                              
defparam Quant_Scan_Matrix_ROM.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                              
defparam Quant_Scan_Matrix_ROM.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                              
defparam Quant_Scan_Matrix_ROM.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Quant_Scan_Matrix_ROM.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// synthesis translate_on
endmodule
  