// 
//  MAC_MPEG2_AV - MPEG-2 hardware implementation for Xilinx multimedia board 
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MPEG2_AV
// 
// MAC_MPEG2_AV is distributed in the hope that it will be useful for further 
// research, but WITHOUT ANY WARRANTY; without even the implied warranty of 
//	MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. MAC_MPEG2_AV is free; you 
// can redistribute it and/or modify it provided that proper reference is provided 
// to the authors. See the documents included in the "doc" folder for further details.
//
//==============================================================================

`include "defines.v"
module Const_ROM_Sample_RAM(
   clock,

   ROM_Enable_I,
   ROM_Address_I,
   ROM_Data_O,

	RAM_Address_I,
	RAM_Data_O,
	RAM_Wen_I,
	RAM_Data_I
);

input 				clock;

input					ROM_Enable_I;
input 	[9:0]		ROM_Address_I;
output 	[15:0]	ROM_Data_O;

input 	[9:0]		RAM_Address_I;
output 	[15:0]	RAM_Data_O;
input 				RAM_Wen_I;
input 	[15:0]	RAM_Data_I;

RAMB16_S18_S18 ROM_RAM_BRAM (
   .DOA(ROM_Data_O),
   .DOB(RAM_Data_O),
   .DOPA(),
   .DOPB(),
   .ADDRA(ROM_Address_I),
   .ADDRB(RAM_Address_I),
   .CLKA(clock),
   .CLKB(clock),
   .DIA(16'h0000),
   .DIB(RAM_Data_I),
   .DIPA(2'b00),
   .DIPB(2'b00),
   .ENA(ROM_Enable_I),
   .ENB(1'b1),
   .SSRA(1'b0),
   .SSRB(1'b0),
   .WEA(1'b0),
   .WEB(RAM_Wen_I)
);

// synthesis attribute WRITE_MODE_B of ROM_RAM_BRAM is "READ_FIRST"

// synthesis attribute INIT_00 of ROM_RAM_BRAM is "256'hffff000000000000000000000000000000000000000000000000000000004947"
// synthesis attribute INIT_01 of ROM_RAM_BRAM is "256'hfffafffafffbfffcfffcfffcfffdfffdfffefffefffeffffffffffffffffffff"
// synthesis attribute INIT_02 of ROM_RAM_BRAM is "256'hffe8ffeaffebffedffeeffeffff1fff2fff3fff4fff5fff6fff7fff8fff9fff9"
// synthesis attribute INIT_03 of ROM_RAM_BRAM is "256'hffcdffceffcfffd1ffd3ffd4ffd6ffd8ffdaffdcffdeffe0ffe1ffe3ffe5ffe7"
// synthesis attribute INIT_04 of ROM_RAM_BRAM is "256'h0028002c002f0032003300350037003800380039003900380038003700360035"
// synthesis attribute INIT_05 of ROM_RAM_BRAM is "256'hff9cffaaffb7ffc3ffcfffdaffe5ffeefff800000007000e0014001a001f0024"
// synthesis attribute INIT_06 of ROM_RAM_BRAM is "256'hfe8afe9bfeadfec0fed2fee4fef6ff09ff1bff2dff3eff4fff5fff6fff7fff8e"
// synthesis attribute INIT_07 of ROM_RAM_BRAM is "256'hfdfdfdf9fdf7fdf7fdfafdfefe05fe0cfe16fe21fe2dfe3afe49fe58fe68fe79"

// synthesis attribute INIT_08 of ROM_RAM_BRAM is "256'h002e0064009700c600f2011a01400161017f019a01b201c701d901e701f301fd"
// synthesis attribute INIT_09 of ROM_RAM_BRAM is "256'hfb54fbaefc09fc62fcbbfd12fd67fdbafe0bfe5afea6feefff35ff78ffb9fff5"
// synthesis attribute INIT_0A of ROM_RAM_BRAM is "256'hf6a4f6cef700f737f774f7b6f7fcf847f895f8e7f93bf991f9e9fa43fa9dfaf8"
// synthesis attribute INIT_0B of ROM_RAM_BRAM is "256'hf909f88bf81af7b5f75ff714f6d5f6a2f67bf65ff64df645f647f652f665f681"
// synthesis attribute INIT_0C of ROM_RAM_BRAM is "256'hf7a9f904fa52fb93fcc7fdeeff070011010e01fd02dd03af0474052a05d1066b"
// synthesis attribute INIT_0D of ROM_RAM_BRAM is "256'hdd33df01e0cee299e460e624e7e3e99ceb4fecfbee9ff03af1ccf354f4d1f643"
// synthesis attribute INIT_0E of ROM_RAM_BRAM is "256'hc2c9c426c591c709c88eca1ecbb9cd5dcf0ad0bfd27ad43bd601d7cbd996db64"
// synthesis attribute INIT_0F of ROM_RAM_BRAM is "256'hb6c5b6e7b71fb76eb7d4b84fb8e0b986ba41bb11bbf5bcecbdf5bf11c03ec17c"

// synthesis attribute INIT_10 of ROM_RAM_BRAM is "256'h0400050A065908000A140CB21000142819652000285132CB400050A265978000"
// synthesis attribute INIT_11 of ROM_RAM_BRAM is "256'h0019002000280032004000500065008000A100CB01000142019602000285032C"
// synthesis attribute INIT_12 of ROM_RAM_BRAM is "256'h000000000001000100010002000200030004000500060008000A000C00100014"
// synthesis attribute INIT_13 of ROM_RAM_BRAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_14 of ROM_RAM_BRAM is "256'h000200040008001000200040008001010204041008421111C71C249299995555"
// synthesis attribute INIT_15 of ROM_RAM_BRAM is "256'h0001000200030008001000200040008001000200040008001000200040000001"
// synthesis attribute INIT_16 of ROM_RAM_BRAM is "256'hbdaec5e4cd9fd4dbdb94e1c5e76bec83f109f4faf853fb14fd3afec4ffb1ffff"
// synthesis attribute INIT_17 of ROM_RAM_BRAM is "256'h0c8f1917259031f13e334a50563e61f76d7478ad839c8e39987fa267abebb504"

// synthesis attribute INIT_18 of ROM_RAM_BRAM is "256'hDA987654321F0E01DCBA987654321001DCBA987654321001DCBA987654321001"
// synthesis attribute INIT_19 of ROM_RAM_BRAM is "256'hDA987654321F0E01DA987654321F0E01DA987654321F0E01DA987654321F0E01"
// synthesis attribute INIT_1A of ROM_RAM_BRAM is "256'hD21F0E02D21F0E02DA987654321F0E01DA987654321F0E01DA987654321F0E01"
// synthesis attribute INIT_1B of ROM_RAM_BRAM is "256'hD21F0E02D21F0E02D21F0E02D21F0E02D21F0E02D21F0E02D21F0E02D21F0E02"
// synthesis attribute INIT_1C of ROM_RAM_BRAM is "256'hFE01CBA987654321FE01DE03DE03DE03DE03DE03DE03DE03D21F0E02D21F0E02"
// synthesis attribute INIT_1D of ROM_RAM_BRAM is "256'hFE024321FE024321FE024321FE024321FE024321FE024321FE02CBA987654321"
// synthesis attribute INIT_1E of ROM_RAM_BRAM is "256'h0E01BA987654321F0E01BA987654321F0E014321FE024321FE024321FE024321"
// synthesis attribute INIT_1F of ROM_RAM_BRAM is "256'hFE024321FE024321FE024321FE024321FE02BA987654321F0E01BA987654321F"
                                                                                                                     
// synthesis attribute INIT_20 of ROM_RAM_BRAM is "256'hFE03FE03FE03FE03FE03FE03FE03FE03FE03FE03FE034321FE024321FE024321"  
// synthesis attribute INIT_21 of ROM_RAM_BRAM is "256'h00000000000000000000000000000000FE03FE03FE03FE03FE03FE03FE03FE03"
// synthesis attribute INIT_22 of ROM_RAM_BRAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_23 of ROM_RAM_BRAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_24 of ROM_RAM_BRAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_25 of ROM_RAM_BRAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_26 of ROM_RAM_BRAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_27 of ROM_RAM_BRAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"

// synthesis translate_off 

defparam ROM_RAM_BRAM.WRITE_MODE_B = "READ_FIRST";

defparam ROM_RAM_BRAM.INIT_00 = 256'hffff000000000000000000000000000000000000000000000000000000004947;
defparam ROM_RAM_BRAM.INIT_01 = 256'hfffafffafffbfffcfffcfffcfffdfffdfffefffefffeffffffffffffffffffff;
defparam ROM_RAM_BRAM.INIT_02 = 256'hffe8ffeaffebffedffeeffeffff1fff2fff3fff4fff5fff6fff7fff8fff9fff9;
defparam ROM_RAM_BRAM.INIT_03 = 256'hffcdffceffcfffd1ffd3ffd4ffd6ffd8ffdaffdcffdeffe0ffe1ffe3ffe5ffe7;
defparam ROM_RAM_BRAM.INIT_04 = 256'h0028002c002f0032003300350037003800380039003900380038003700360035;
defparam ROM_RAM_BRAM.INIT_05 = 256'hff9cffaaffb7ffc3ffcfffdaffe5ffeefff800000007000e0014001a001f0024;
defparam ROM_RAM_BRAM.INIT_06 = 256'hfe8afe9bfeadfec0fed2fee4fef6ff09ff1bff2dff3eff4fff5fff6fff7fff8e;
defparam ROM_RAM_BRAM.INIT_07 = 256'hfdfdfdf9fdf7fdf7fdfafdfefe05fe0cfe16fe21fe2dfe3afe49fe58fe68fe79;

defparam ROM_RAM_BRAM.INIT_08 = 256'h002e0064009700c600f2011a01400161017f019a01b201c701d901e701f301fd;
defparam ROM_RAM_BRAM.INIT_09 = 256'hfb54fbaefc09fc62fcbbfd12fd67fdbafe0bfe5afea6feefff35ff78ffb9fff5;
defparam ROM_RAM_BRAM.INIT_0A = 256'hf6a4f6cef700f737f774f7b6f7fcf847f895f8e7f93bf991f9e9fa43fa9dfaf8;
defparam ROM_RAM_BRAM.INIT_0B = 256'hf909f88bf81af7b5f75ff714f6d5f6a2f67bf65ff64df645f647f652f665f681;
defparam ROM_RAM_BRAM.INIT_0C = 256'hf7a9f904fa52fb93fcc7fdeeff070011010e01fd02dd03af0474052a05d1066b;
defparam ROM_RAM_BRAM.INIT_0D = 256'hdd33df01e0cee299e460e624e7e3e99ceb4fecfbee9ff03af1ccf354f4d1f643;
defparam ROM_RAM_BRAM.INIT_0E = 256'hc2c9c426c591c709c88eca1ecbb9cd5dcf0ad0bfd27ad43bd601d7cbd996db64;
defparam ROM_RAM_BRAM.INIT_0F = 256'hb6c5b6e7b71fb76eb7d4b84fb8e0b986ba41bb11bbf5bcecbdf5bf11c03ec17c;

defparam ROM_RAM_BRAM.INIT_10 = 256'h0400050A065908000A140CB21000142819652000285132CB400050A265978000;
defparam ROM_RAM_BRAM.INIT_11 = 256'h0019002000280032004000500065008000A100CB01000142019602000285032C;
defparam ROM_RAM_BRAM.INIT_12 = 256'h000000000001000100010002000200030004000500060008000A000C00100014;
defparam ROM_RAM_BRAM.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ROM_RAM_BRAM.INIT_14 = 256'h000200040008001000200040008001010204041008421111C71C249299995555;
defparam ROM_RAM_BRAM.INIT_15 = 256'h0001000200030008001000200040008001000200040008001000200040000001;
defparam ROM_RAM_BRAM.INIT_16 = 256'hbdaec5e4cd9fd4dbdb94e1c5e76bec83f109f4faf853fb14fd3afec4ffb1ffff;
defparam ROM_RAM_BRAM.INIT_17 = 256'h0c8f1917259031f13e334a50563e61f76d7478ad839c8e39987fa267abebb504;
                                                                                                  
defparam ROM_RAM_BRAM.INIT_18 = 256'hDA987654321F0E01DCBA987654321001DCBA987654321001DCBA987654321001;
defparam ROM_RAM_BRAM.INIT_19 = 256'hDA987654321F0E01DA987654321F0E01DA987654321F0E01DA987654321F0E01;
defparam ROM_RAM_BRAM.INIT_1A = 256'hD21F0E02D21F0E02DA987654321F0E01DA987654321F0E01DA987654321F0E01;
defparam ROM_RAM_BRAM.INIT_1B = 256'hD21F0E02D21F0E02D21F0E02D21F0E02D21F0E02D21F0E02D21F0E02D21F0E02;
defparam ROM_RAM_BRAM.INIT_1C = 256'hFE01CBA987654321FE01DE03DE03DE03DE03DE03DE03DE03D21F0E02D21F0E02;
defparam ROM_RAM_BRAM.INIT_1D = 256'hFE024321FE024321FE024321FE024321FE024321FE024321FE02CBA987654321;
defparam ROM_RAM_BRAM.INIT_1E = 256'h0E01BA987654321F0E01BA987654321F0E014321FE024321FE024321FE024321;
defparam ROM_RAM_BRAM.INIT_1F = 256'hFE024321FE024321FE024321FE024321FE02BA987654321F0E01BA987654321F;
                          
defparam ROM_RAM_BRAM.INIT_20 = 256'hFE03FE03FE03FE03FE03FE03FE03FE03FE03FE03FE034321FE024321FE024321;
defparam ROM_RAM_BRAM.INIT_21 = 256'h00000000000000000000000000000000FE03FE03FE03FE03FE03FE03FE03FE03;
defparam ROM_RAM_BRAM.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ROM_RAM_BRAM.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ROM_RAM_BRAM.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ROM_RAM_BRAM.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ROM_RAM_BRAM.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam ROM_RAM_BRAM.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                     
// synthesis translate_on

endmodule
