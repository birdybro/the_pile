// 
//  MAC_MPEG2_AV - MPEG-2 hardware implementation for Xilinx multimedia board 
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MPEG2_AV
// 
// MAC_MPEG2_AV is distributed in the hope that it will be useful for further 
// research, but WITHOUT ANY WARRANTY; without even the implied warranty of 
//	MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. MAC_MPEG2_AV is free; you 
// can redistribute it and/or modify it provided that proper reference is provided 
// to the authors. See the documents included in the "doc" folder for further details.
//
//==============================================================================

`include "defines.v"
module bram(clock, wren_a, wren_b, address_a, address_b, data_in_a, data_in_b, data_out_a, data_out_b);

input clock;
input wren_a, wren_b;
input [`IDCT_ADDR_WIDTH-1:0] address_a, address_b;
input [`IDCT_DATA_WIDTH-1:0] data_in_a, data_in_b;
output [`IDCT_DATA_WIDTH-1:0] data_out_a, data_out_b;

wire [31:0] dummy_a, dummy_b;

assign data_out_a = dummy_a[`IDCT_DATA_WIDTH-1:0];
assign data_out_b = dummy_b[`IDCT_DATA_WIDTH-1:0];

// Instantiate the RAM
RAMB16_S36_S36 instance_bram (
      .DOA(dummy_a),     
      .DOB(dummy_b),     
      .DOPA(),		   		 
      .DOPB(),					
      .ADDRA({2'b00,address_a}),
      .ADDRB({2'b00,address_b}),
      .CLKA(clock),  
      .CLKB(clock),  
      .DIA({8'h00,data_in_a}),    
      .DIB({8'h00,data_in_b}),    
      .DIPA(4'h0),  
      .DIPB(4'h0),  
      .ENA(1'b1),
      .ENB(1'b1),
      .SSRA(1'b0),  
      .SSRB(1'b0),  
      .WEA(wren_a),    
      .WEB(wren_b)     
   );

// synthesis attribute INIT_00 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_01 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_02 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_03 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_04 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_05 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_06 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_07 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_08 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_09 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0A of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0B of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0C of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0D of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0E of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0F of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_10 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_11 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_12 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_13 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_14 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_15 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_16 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_17 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_18 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_19 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1A of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1B of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1C of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1D of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1E of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1F of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_20 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_21 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_22 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_23 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_24 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_25 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_26 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_27 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_28 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_29 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2A of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2B of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2C of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2D of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2E of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2F of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_30 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_31 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_32 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_33 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_34 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_35 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_36 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_37 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_38 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_39 of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3A of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3B of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3C of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3D of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3E of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3F of instance_bram is "256'h0000000000000000000000000000000000000000000000000000000000000000"

// synthesis translate_off
/*
defparam instance_bram.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam instance_bram.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
*/
// synthesis translate_on

endmodule
