// 
//  MAC_MPEG2_AV - MPEG-2 hardware implementation for Xilinx multimedia board 
//  Copyright (C) 2007 McMaster University
// 
//==============================================================================
// 
// This file is part of MAC_MPEG2_AV
// 
// MAC_MPEG2_AV is distributed in the hope that it will be useful for further 
// research, but WITHOUT ANY WARRANTY; without even the implied warranty of 
//	MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. MAC_MPEG2_AV is free; you 
// can redistribute it and/or modify it provided that proper reference is provided 
// to the authors. See the documents included in the "doc" folder for further details.
//
//==============================================================================

`include "defines.v"
module MC_Prediction_Buffer(
   clock,
   Write_En_A_I,
   Address_A_I,
   Data_A_I,
   Data_A_O,
   Write_En_B_I,
   Address_B_I,
   Data_B_I,
   Data_B_O
);

input             clock;
input             Write_En_A_I;
input    [9:0]    Address_A_I;
input    [15:0]   Data_A_I;
output   [15:0]   Data_A_O;
input             Write_En_B_I;
input    [9:0]    Address_B_I;
input    [15:0]   Data_B_I;
output   [15:0]   Data_B_O;

RAMB16_S18_S18 Buffer_RAM (
   .DOA(Data_A_O),
   .DOB(Data_B_O),
   .DOPA(),
   .DOPB(),
   .ADDRA(Address_A_I),
   .ADDRB(Address_B_I),
   .CLKA(clock),
   .CLKB(clock),
   .DIA(Data_A_I),
   .DIB(Data_B_I),
   .DIPA(2'b00),
   .DIPB(2'b00),
   .ENA(1'b1),
   .ENB(1'b1),
   .SSRA(1'b0),
   .SSRB(1'b0),
   .WEA(Write_En_A_I),
   .WEB(Write_En_B_I)
);
  
// synthesis attribute INIT_00 of Buffer_RAM is "256'h8D8C8B8A8988100F0E0D0C0B870A858611120809848306078205030481800102"
// synthesis attribute INIT_01 of Buffer_RAM is "256'h9C9B9A9921201F1E22231D1C1A1B979695949819181793929190151614138F8E"
// synthesis attribute INIT_02 of Buffer_RAM is "256'hACABAAA931302F2EA8A7A6A5A4A3A2A12B2A29282D2C272632332524A09F9E9D"
// synthesis attribute INIT_03 of Buffer_RAM is "256'hBCBBBAB941403F3EB8B7B6B5B4B3B2B13B3A39383D3C373642433534B0AFAEAD"
// synthesis attribute INIT_04 of Buffer_RAM is "256'hCCCBCAC951504F4EC8C7C6C5C4C3C2C14B4A49484D4C474652534544C0BFBEBD"
// synthesis attribute INIT_05 of Buffer_RAM is "256'hDCDBDAD961605F5ED8D7D6D5D4D3D2D15B5A59585D5C575662ff5554D0CFCECD"
// synthesis attribute INIT_06 of Buffer_RAM is "256'hEEEDECEBEAE9706F6E6DE8E7E6E5E4E3E2E16A6968676C6B66656463E0DFDEDD"
// synthesis attribute INIT_07 of Buffer_RAM is "256'h8B8A0E890D880C870B860A85098408830782818083800804828106050302F0EF"
                                                                                                                     
// synthesis attribute INIT_08 of Buffer_RAM is "256'h0A010005010303020B010C0100060D0100030401030102010002010100014000"  
// synthesis attribute INIT_09 of Buffer_RAM is "256'h0E010F0101040203000705021001410008010004090102020501010206010701"
// synthesis attribute INIT_0A of Buffer_RAM is "256'h06020008030301051201130100091401150107020204000A04030802000B0402"
// synthesis attribute INIT_0B of Buffer_RAM is "256'h1701180119011A01000C000D000E000F0106010702050304050309020A021101"
// synthesis attribute INIT_0C of Buffer_RAM is "256'h001100120013001400150016001700180019001A001B001C001D001E001F1601"
// synthesis attribute INIT_0D of Buffer_RAM is "256'h0109010A010B010C010D010E0020002100220023002400250026002700280010"
// synthesis attribute INIT_0E of Buffer_RAM is "256'h1C011D011E011F010B020C020D020E020F0210020603010F0110011101120108"
// synthesis attribute INIT_0F of Buffer_RAM is "256'h000000000000000091FF9A96090A819E07088A880506868403048E8C01021B01"
                                                                                                                     
// synthesis attribute INIT_10 of Buffer_RAM is "256'h8E8D8C8B8A890F0E0D88878685840C0B0A090807838206050481101103800102"
// synthesis attribute INIT_11 of Buffer_RAM is "256'h222321209A999897969594931D1C1B1A19189C9B92171E1F161591901314128F"
// synthesis attribute INIT_12 of Buffer_RAM is "256'h373631303C3D2F2EAAA9A82BA7A62C2D2A292728A4A3A2A1A5262524A09F9E9D"
// synthesis attribute INIT_13 of Buffer_RAM is "256'h474641404B4C3F3EB4B3ffB2ffB1B0ff3B3A3938AFAEADffffACABff35343332"
// synthesis attribute INIT_14 of Buffer_RAM is "256'h52515655504F5B5C4E4DC0BFBEBDBCff4A4948ffffBBBAB9B8B7B6B545444342"
// synthesis attribute INIT_15 of Buffer_RAM is "256'h62616665605F6Bff5E5DD0CFCECDCCCBCAC95A595857C8C7C6C5C4C3C2C15453"
// synthesis attribute INIT_16 of Buffer_RAM is "256'h7372717075746F6E6D6CE0DFDEDDDCDBDAD96A696867D8D7D6D5D4D3D2D16463"
// synthesis attribute INIT_17 of Buffer_RAM is "256'h000000000000000091FF8101F0EFEEEDECEBEAE979787776E8E7E6E5E4E3E2E1"
                                                                                                                     
// synthesis attribute INIT_18 of Buffer_RAM is "256'h0101000F000E04020203000D000C000900080A01010309010005000400020001"
// synthesis attribute INIT_19 of Buffer_RAM is "256'h04010006000703010102010403020C010D01000A000B0B010105020100034000"
// synthesis attribute INIT_1A of Buffer_RAM is "256'h14011501070204030802100102040F010E010502410002020601080107010501"
// synthesis attribute INIT_1B of Buffer_RAM is "256'h1701180119011A010106010702050304050309020A0211010602030312011301"
// synthesis attribute INIT_1C of Buffer_RAM is "256'h001100120013001400150016001700180019001A001B001C001D001E001F1601"
// synthesis attribute INIT_1D of Buffer_RAM is "256'h0109010A010B010C010D010E0020002100220023002400250026002700280010"
// synthesis attribute INIT_1E of Buffer_RAM is "256'h1C011D011E011F010B020C020D020E020F0210020603010F0110011101120108"
// synthesis attribute INIT_1F of Buffer_RAM is "256'h0809868706078485040582830203810191FF9206819A0405880382028A011B01"
                                                                                                                     
// synthesis attribute INIT_20 of Buffer_RAM is "256'h18199495929390911617141512138E8F1A1B10118C8D8A8B0C0D88890E0F0A0B"
// synthesis attribute INIT_21 of Buffer_RAM is "256'h81028001ffE1ff25ff24A0A19E9F9C9D9A9B21221F201D1E23ff1Cff98999697"
// synthesis attribute INIT_22 of Buffer_RAM is "256'h8F908D8E10110F0F8B8C8A0D88890B0C0E0E870A858608098407050683048203"
// synthesis attribute INIT_23 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_24 of Buffer_RAM is "256'hB4B89CAC10110E0F12130C0D94A88CB0080990A084880607BC050A0B03040102"
// synthesis attribute INIT_25 of Buffer_RAM is "256'h2E2F202192A2868A91A185891C1D1A1B83BF98A4181916171E1F141582BE81BD"
// synthesis attribute INIT_26 of Buffer_RAM is "256'h3637303197AB8FB396AA8EB22C2D2A2B95A98DB193A3878B2627242528292223"
// synthesis attribute INIT_27 of Buffer_RAM is "256'h80809BA7B7BB9FAF3E3F3C3DB6BA9EAE3A3B3839B5B99DAD9AA699A534353233"
                                                                                                                     
// synthesis attribute INIT_28 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_29 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2A of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2B of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2C of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2D of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2E of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2F of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
                                                                                                                     
// synthesis attribute INIT_30 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_31 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_32 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_33 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_34 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_35 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_36 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_37 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
                                                                                                                     
// synthesis attribute INIT_38 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_39 of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3A of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3B of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3C of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3D of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3E of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3F of Buffer_RAM is "256'h0000000000000000000000000000000000000000000000000000000000000000"

// synthesis translate_off 
 
defparam Buffer_RAM.INIT_00 = 256'h8D8C8B8A8988100F0E0D0C0B870A858611120809848306078205030481800102;
defparam Buffer_RAM.INIT_01 = 256'h9C9B9A9921201F1E22231D1C1A1B979695949819181793929190151614138F8E;
defparam Buffer_RAM.INIT_02 = 256'hACABAAA931302F2EA8A7A6A5A4A3A2A12B2A29282D2C272632332524A09F9E9D;
defparam Buffer_RAM.INIT_03 = 256'hBCBBBAB941403F3EB8B7B6B5B4B3B2B13B3A39383D3C373642433534B0AFAEAD;
defparam Buffer_RAM.INIT_04 = 256'hCCCBCAC951504F4EC8C7C6C5C4C3C2C14B4A49484D4C474652534544C0BFBEBD;
defparam Buffer_RAM.INIT_05 = 256'hDCDBDAD961605F5ED8D7D6D5D4D3D2D15B5A59585D5C575662ff5554D0CFCECD;
defparam Buffer_RAM.INIT_06 = 256'hEEEDECEBEAE9706F6E6DE8E7E6E5E4E3E2E16A6968676C6B66656463E0DFDEDD;
defparam Buffer_RAM.INIT_07 = 256'h8B8A0E890D880C870B860A85098408830782818083800804828106050302F0EF;
                                                                                                                                         
defparam Buffer_RAM.INIT_08 = 256'h0A010005010303020B010C0100060D0100030401030102010002010100014000;
defparam Buffer_RAM.INIT_09 = 256'h0E010F0101040203000705021001410008010004090102020501010206010701;
defparam Buffer_RAM.INIT_0A = 256'h06020008030301051201130100091401150107020204000A04030802000B0402;
defparam Buffer_RAM.INIT_0B = 256'h1701180119011A01000C000D000E000F0106010702050304050309020A021101;
defparam Buffer_RAM.INIT_0C = 256'h001100120013001400150016001700180019001A001B001C001D001E001F1601;
defparam Buffer_RAM.INIT_0D = 256'h0109010A010B010C010D010E0020002100220023002400250026002700280010;
defparam Buffer_RAM.INIT_0E = 256'h1C011D011E011F010B020C020D020E020F0210020603010F0110011101120108;
defparam Buffer_RAM.INIT_0F = 256'h000000000000000091FF9A96090A819E07088A880506868403048E8C01021B01;

defparam Buffer_RAM.INIT_10 = 256'h8E8D8C8B8A890F0E0D88878685840C0B0A090807838206050481101103800102;
defparam Buffer_RAM.INIT_11 = 256'h222321209A999897969594931D1C1B1A19189C9B92171E1F161591901314128F;
defparam Buffer_RAM.INIT_12 = 256'h373631303C3D2F2EAAA9A82BA7A62C2D2A292728A4A3A2A1A5262524A09F9E9D;
defparam Buffer_RAM.INIT_13 = 256'h474641404B4C3F3EB4B3ffB2ffB1B0ff3B3A3938AFAEADffffACABff35343332;
defparam Buffer_RAM.INIT_14 = 256'h52515655504F5B5C4E4DC0BFBEBDBCff4A4948ffffBBBAB9B8B7B6B545444342;
defparam Buffer_RAM.INIT_15 = 256'h62616665605F6Bff5E5DD0CFCECDCCCBCAC95A595857C8C7C6C5C4C3C2C15453;
defparam Buffer_RAM.INIT_16 = 256'h7372717075746F6E6D6CE0DFDEDDDCDBDAD96A696867D8D7D6D5D4D3D2D16463;
defparam Buffer_RAM.INIT_17 = 256'h000000000000000091FF8101F0EFEEEDECEBEAE979787776E8E7E6E5E4E3E2E1;

defparam Buffer_RAM.INIT_18 = 256'h0101000F000E04020203000D000C000900080A01010309010005000400020001;
defparam Buffer_RAM.INIT_19 = 256'h04010006000703010102010403020C010D01000A000B0B010105020100034000;
defparam Buffer_RAM.INIT_1A = 256'h14011501070204030802100102040F010E010502410002020601080107010501;
defparam Buffer_RAM.INIT_1B = 256'h1701180119011A010106010702050304050309020A0211010602030312011301;
defparam Buffer_RAM.INIT_1C = 256'h001100120013001400150016001700180019001A001B001C001D001E001F1601;
defparam Buffer_RAM.INIT_1D = 256'h0109010A010B010C010D010E0020002100220023002400250026002700280010;
defparam Buffer_RAM.INIT_1E = 256'h1C011D011E011F010B020C020D020E020F0210020603010F0110011101120108;
defparam Buffer_RAM.INIT_1F = 256'h0809868706078485040582830203810191FF9206819A0405880382028A011B01;

defparam Buffer_RAM.INIT_20 = 256'h18199495929390911617141512138E8F1A1B10118C8D8A8B0C0D88890E0F0A0B;
defparam Buffer_RAM.INIT_21 = 256'h81028001ffE1ff25ff24A0A19E9F9C9D9A9B21221F201D1E23ff1Cff98999697;
defparam Buffer_RAM.INIT_22 = 256'h8F908D8E10110F0F8B8C8A0D88890B0C0E0E870A858608098407050683048203;
defparam Buffer_RAM.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_24 = 256'hB4B89CAC10110E0F12130C0D94A88CB0080990A084880607BC050A0B03040102;
defparam Buffer_RAM.INIT_25 = 256'h2E2F202192A2868A91A185891C1D1A1B83BF98A4181916171E1F141582BE81BD;
defparam Buffer_RAM.INIT_26 = 256'h3637303197AB8FB396AA8EB22C2D2A2B95A98DB193A3878B2627242528292223;
defparam Buffer_RAM.INIT_27 = 256'h80809BA7B7BB9FAF3E3F3C3DB6BA9EAE3A3B3839B5B99DAD9AA699A534353233;
                                                                                                  
defparam Buffer_RAM.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                  
defparam Buffer_RAM.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
                                                                                                  
defparam Buffer_RAM.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam Buffer_RAM.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// synthesis translate_on
endmodule
